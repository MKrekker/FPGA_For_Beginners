$date
  Thu Nov 18 15:09:54 2021
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module d_ff $end
$var reg 1 ! d_in $end
$var reg 1 " clk $end
$var reg 1 # q_o $end
$upscope $end
$enddefinitions $end
#0
U!
1"
U#
#5000000000
0"
